// $Id: $
// File name:   bit_stuffer_detect.sv
// Created:     4/29/2020
// Author:      Wang-Ning Lo
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Bit Stuffer Detector
